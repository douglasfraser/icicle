// Defines for Olimex iCE40HX8K-EVB development board
//`define FLASH
